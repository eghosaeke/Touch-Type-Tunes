BZh91AY&SYi��� G߀Px����������P���3�nr�ۡ$���j#`�i�Ѡ ����3J��e=L�F� 21�2 " SB#�̈��  ��hhɉ�	���0 �`�0�$�S���i���  4���$��"�	����ңH7��/p�%f�{]�bV�X|������QW��ɍ��t*�爗��I��VM{��a��P�l�ݷ�A�3�>4�/ДT�jY xJ�A ���f���0�3�<	<�&��K�\�0k@��-w�ݷ���R���n����L�fO6v��Q�ٗfXh���j顖|�N�fC��2z:i�7�g�gEL��t-������`�f�-�ˡJ8�aڊ��-�X���v��x���%�@�S���aC^",�fbf�Ҷ��r���>�1^�R9#���J���dn����Be@O��sTф��2�k�}�wgs�a�2���a8�R}��^�������+���/`�<B-���Yɋ,_��kU��`���VoG������7*HR5j�z�퇺��*q�P
g	Bk(����*d�����a��u*8t�ƑT�5E�ZK	穀� Q��a�� ��0�^��q���;�Z�*���pZ<��e����	�b�C�ï�g�N6��}5�l.��6�.��&!.��9S):� ZL��Ahh���7�.�,Pqj,S����FJl�`��&��j�B`����]a�8[@�}[�E�lɲ�'��n2C�Ĳ��#fW��!��\��7M�)m;��<5�J�Q�:��|�j�Р���-ٍnM22�bA�ٙYU���xb\��1�-Ib��E3I����O]dr0,pp�HT���!Ŗ�u�-�̾��+�,,T��C�]��BA�&3