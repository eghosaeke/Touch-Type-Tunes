BZh91AY&SY���T �_�Px����������P�rT���0��'�B��E4d�@ڏP hCCjѓ �`A��2`�S$#DHSɤި  ���101��&$Ja	���d�O�O�6���a��CܒSBU ���?c�a��h���D�ہ|$�Z0
0<\�cmF���n�|\�ߛu^��G��t��ڦ1Y�sc��-HIM4�ћz��~��f�0�&�QW5Ņ��P���`kƥ�� δ�Ӛ@�0� ����}�.�*�������:qABb�[�F���e�K��YNX꺾;[fYI}T�����H�r3,��mEq�<Ԕ�Tt	��a�j�	���K�2�2-q��������K��)�:�B��I%!1�F��$o�j�И�k#�ک*U������R�LKm
S*��JGB��l��*��f�bH���9����Kh�io˂#ǡ�V�E*B2�dH��?{�}`d���|F��-xl=���&�|&̙���ArE�=�1���#,�
A����U��QV�"gCZ+�"�jq*�"Ũk�jR�4F�a��� ���I9Nt���Zx�e�2�C����N��u�hR��;YĮ���#����PTб���y�@i�}�fE�T�`{���w��,��^B�,[����� �M�$#�ņ�:63=Ć�(u��1Q�2��a+B�)+h����Ϟ��<�:m���:�@����: �Y���)�˸0*m-� h$,%#@2�X��X`0��B��0�!�c��lj`��# �#��`���,<��I�6tڄ�i��n03�#��䦪xm6� �� �^�:npj�>��g���B�a�ϩBA#�ZT�d���c`�I��, ��"C�f�c4�l�gh��9<
LR��*j���	�Lʆb�=����K�@�KS��I��ļZF��^)1y�n$m�5�2�Z��1�m��m���6�����A�a���3�]��BB���P