BZh91AY&SY�y�� �_�Px����������P�v�g*%T�(@�4��ѩ�=#Ѩڍ 4�M��i�I@   �h  ��Q�P4i�F�  �4 挘� ���F	� �$��iM?M2SѨ=OP  ��d3Ԑ��+L��M*�H�����)$���Ͷ ���h0���4�i��v��>K%��d���@#"���IW{���W@����T+Ŵ�8�^�^>8L�7"iW9[P$N� ��M6q�L	��c�.~�h� ���ݡq��"����ܙ!a#KL�ӑ �A�5���i Hr�jZET^B��*�Y V���A �L(a!�1�y���!+@����yI�T�R"(��ĵ @�� 0�&�ͦ���^��J�������EC�҅u"����0'@'��n�Tô;'�7�%`
���[z��J8W���㳅�?�@��R�Y�8|i��IXN�'o[��&5a^���;ױ3�:�M����x�����ؠ��F�y���P�$�ց�%�3�c��b$�?�I�"!�R�b*cc`��+7llD,!F j�zB�V8�Y���2}��J(�&��y��(UgC�3��\QQ6��zf�߈`m7�@��Z+��8��D6!}Ƞ�>c�*=O���X^ሎt����A�Z����D��%��ߴ
�S@`a��Ԭ4�7=/�0�Yc_�N��L�}��
����u�'�*����o�'RA@Ta��9t�t�M��{3*S@!b:*i��*�Ԉje`J	c��� wH��@��w���N\5#���1��+����1ǽ�\�Sk��H	z7�&�!X��sC5࡜k�#�f$z�S>�Q�J����G9g\$cI��eVu���c���Vo�@bIk�{�E�ս�w��եIEK��+��w��392����h�U;��5O�&9TMw���-�W�rE8P��y��